--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   10:59:25 05/19/2020
-- Design Name:   
-- Module Name:   D:/zeta/hopeitsfinal/MULTITEST.vhd
-- Project Name:  hopeitsfinal
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Project_MultiC
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY MULTITEST IS
END MULTITEST;
 
ARCHITECTURE behavior OF MULTITEST IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Project_MultiC
    PORT(
         Clk : IN  std_logic;
         Rst : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal Clk : std_logic := '0';
   signal Rst : std_logic := '0';

   -- Clock period definitions
   constant Clk_period : time := 150 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Project_MultiC PORT MAP (
          Clk => Clk,
          Rst => Rst
        );

   -- Clock process definitions
   Clk_process :process
   begin
		Clk <= '0';
		wait for Clk_period/2;
		Clk <= '1';
		wait for Clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
		Rst <= '1';
		wait for Clk_period*1;
		
		
		Rst <= '0';
		wait for Clk_period*5;
		
      wait;
   end process;

END;
